module ADDW();

endmodule